Simulation 4 - 20 mA

* TL074 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.01 ON 06/16/89 AT 13:08
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TL074    1 2 3 4 5
*
  C1   11 12 3.498E-12
  C2    6  7 15.00E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 4.715E6 -5E6 5E6 5E6 -5E6
  GA    6  0 11 12 282.8E-6
  GCM   0  6 10 99 8.942E-9
  ISS   3 10 DC 195.0E-6
  HLIM 90  0 VLIM 1K
  J1   11  2 10 JX
  J2   12  1 10 JX
  R2    6  9 100.0E3
  RD1   4 11 3.536E3
  RD2   4 12 3.536E3
  RO1   8  5 150
  RO2   7 99 150
  RP    3  4 2.143E3
  RSS  10 99 1.026E6
  VB    9  0 DC 0
  VC    3 53 DC 2.200
  VE   54  4 DC 2.200
  VLIM  7  8 DC 0
  VLP  91  0 DC 25
  VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=15.00E-12 BETA=270.1E-6 VTO=-1)
.ENDS

* 
.MODEL QBC337 NPN( 
+    IS = 4.13E-14 
+    NF = 0.9822 
+    ISE = 3.534E-15 
+    NE = 1.35 
+    BF = 292.4 
+    IKF = 0.9 
+    VAF = 145.7 
+    NR = 0.982 
+    ISC = 1.957E-13 
+    NC = 1.3 
+    BR = 23.68 
+    IKR = 0.1 
+    VAR = 20 
+    RB = 60 
+    IRB = 0.0002 
+    RBM = 8 
+    RE = 0.1129 
+    RC = 0.25 
+    XTB = 0 
+    EG = 1.11 
+    XTI = 3 
+    CJE = 3.799E-11 
+    VJE = 0.6752 
+    MJE = 0.3488 
+    TF = 5.4E-10 
+    XTF = 4 
+    VTF = 4.448 
+    ITF = 0.665 
+    PTF = 90 
+    CJC = 1.355E-11 
+    VJC = 0.3523 
+    MJC = 0.3831 
+    XCJC = 0.455 
+    TR = 3E-08 
+    CJS = 0 
+    VJS = 0.75 
+    MJS = 0.333 
+    FC = 0.643)
*

**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*    Modeling services provided by   *
* Interface Technologies www.i-t.com *
**************************************
.MODEL bd136 pnp
+IS=1e-09 BF=681.414 NF=0.85 VAF=10
+IKF=0.196957 ISE=1e-08 NE=1.57381 BR=56.5761
+NR=1.5 VAR=0.975138 IKR=0.952908 ISC=1e-08
+NC=3.58666 RB=40.4245 IRB=0.1 RBM=0.106663
+RE=0.00034585 RC=1.31191 XTB=22.4074 XTI=1
+EG=1.05 CJE=1e-11 VJE=0.75 MJE=0.33
+TF=1e-09 XTF=1 VTF=10 ITF=0.01
+CJC=1e-11 VJC=0.75 MJC=0.33 XCJC=0.9
+FC=0.5 CJS=0 VJS=0.75 MJS=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
* Model generated on Feb 22, 2004
* Model format: SPICE3

V24 2 0 DC 24
VM5  1 0 DC -5
VZ 10 11 DC 0

XOP 3 4 2 1 5 TL074

R1 6 0 150
R2 4 6 10k
R3 7 2 820
R4 2 9 43
R5 11 6 100
R6 8 0 2200

*C1 1 5 100p

Q1 7 5 8 QBC337
Q2 10 7 9 bd136

VC 3 0 3

.dc VC .6 3 .01

.control
run
plot v(5)
plot VZ#branch
print VZ#branch
.endc
.end
